module float_add_